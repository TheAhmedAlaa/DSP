module main (
    A,B,C,D,clk,carryin,opmode_b,BCIN,RSTA,RSTB,RSTM,RSTP,RSTC,RSTD,RSTCARRYIN,RSTOPMODE,
    CEA,CEB,CEM,CEP,CEC,CED,CECARRYIN,CEOPMODE,PCIN,BCOUT,PCOUT,P,M,CARRYOUT,CARRYOUTF
);
input [17:0] A,B,D,BCIN;
input [47:0] C,PCIN;
input [7:0] opmode_b;
input clk,carryin,RSTA,RSTB,RSTM,RSTP,RSTC,RSTD,RSTCARRYIN,RSTOPMODE,CEA,CEB,CEM,CEP,CEC,CED,CECARRYIN,CEOPMODE;
output [17:0] BCOUT;
output [47:0] PCOUT,P;
output [35:0] M; 
output CARRYOUT,CARRYOUTF;
parameter A0REG=0;
parameter A1REG=1;
parameter B0REG=0;
parameter B1REG=1;
parameter CREG=1;
parameter DREG=1;
parameter MREG=1;
parameter PREG=1;
parameter CARRYINREG=1; 
parameter CARRYOUTREG=1;
parameter OPMODEREG=1;
parameter CARRYINSEL="OPMODE5";
parameter B_INPUT="DIRECT";
parameter RSTTYPE="SYNC";
wire [17:0] B1,B0,D1,A1;
wire [47:0] C1;
wire [17:0]AS,B1a,ACOUT; 
wire [47:0] D_A_B;
wire [47:0]XOUT,ZOUT;
wire [7:0] opmode;
wire [47:0] zero=48'd0;
wire CYO;
wire [47:0] P__REG;
wire CIN_O;
wire CIN_CIN;
wire [35:0]multiply;
wire [17:0] addd,subb;
block #(.Width(8),.RSTTYPE(RSTTYPE)) OPMODE_REG(.in(opmode_b),.clk(clk),.rst(RSTOPMODE),.ce(CEOPMODE),.sel(OPMODEREG),.out(opmode));
mux_B #(.Width(18),.B_INPUT(B_INPUT)) B_BCIN(.in0(B),.in1(BCIN),.out(B0));
block #(.Width(18),.RSTTYPE(RSTTYPE)) D_REG(.in(D),.clk(clk),.rst(RSTD),.ce(CED),.sel(DREG),.out(D1));
block #(.Width(18),.RSTTYPE(RSTTYPE)) B0_REG(.in(B0),.clk(clk),.rst(RSTB),.ce(CEB),.sel(B0REG),.out(B1));
block #(.Width(18),.RSTTYPE(RSTTYPE)) A0_REG(.in(A),.clk(clk),.rst(RSTA),.ce(CEA),.sel(A0REG),.out(A1));
block #(.Width(48),.RSTTYPE(RSTTYPE)) C_REG(.in(C),.clk(clk),.rst(RSTC),.ce(CEC),.sel(CREG),.out(C1));
assign addd=D1+B1;
assign subb=D1-B1;
mux #(.Width(18)) ADDER_SUB(.in0(addd),.in1(subb),.sel(opmode[6]),.out(AS));
mux #(.Width(18)) opmode4(.in0(B1),.in1(AS),.sel(opmode[4]),.out(B1a));
block #(.Width(18),.RSTTYPE(RSTTYPE)) B1_REG(.in(B1a),.clk(clk),.rst(RSTB),.ce(CEB),.sel(B1REG),.out(BCOUT));
block #(.Width(18),.RSTTYPE(RSTTYPE)) A1_REG(.in(A1),.clk(clk),.rst(RSTA),.ce(CEA),.sel(A1REG),.out(ACOUT));
assign multiply = ACOUT * BCOUT;
block #(.Width(36),.RSTTYPE(RSTTYPE)) M_REG(.in(multiply),.clk(clk),.rst(RSTM),.ce(CEM),.sel(MREG),.out(M));
assign D_A_B={D1[11:0],ACOUT[17:0],BCOUT[17:0]};
mux_4 #(.Width(48)) X(.in0(zero),.in1({12'b0,M}),.in2(PCOUT),.in3(D_A_B),.sel(opmode[1:0]),.out(XOUT));
mux_4 #(.Width(48)) Z(.in0(zero),.in1(PCIN),.in2(PCOUT),.in3(C1),.sel(opmode[3:2]),.out(ZOUT));
mux_CI #(.Width(1),.CARRYINSEL(CARRYINSEL)) CARRY_CASCADE(.in0(carryin),.in1(opmode[5]),.out(CIN_O));
block #(.Width(1),.RSTTYPE(RSTTYPE)) CYI(.in(CIN_O),.clk(clk),.rst(RSTCARRYIN),.ce(CECARRYIN),.sel(CARRYINREG),.out(CIN_CIN));
ADDITION ADD (.XOUT(XOUT),.ZOUT(ZOUT),.opmode7(opmode[7]),.CIN(CIN_CIN),.CYO(CYO),.P(P__REG));
block #(.Width(1),.RSTTYPE(RSTTYPE)) CYO_(.in(CYO),.clk(clk),.rst(RSTCARRYIN),.ce(CECARRYIN),.sel(CARRYOUTREG),.out(CARRYOUT));
assign CARRYOUTF=CARRYOUT;
block #(.Width(48),.RSTTYPE(RSTTYPE)) P_REG(.in(P__REG),.clk(clk),.rst(RSTP),.ce(CEP),.sel(PREG),.out(P));
assign PCOUT=P;
endmodule 